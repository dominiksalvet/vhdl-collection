-- Still under developing!
