-- Still under development!
